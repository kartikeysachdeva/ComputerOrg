module top (CLOCK_50, SW, KEY, LEDR);

    input CLOCK_50;             // DE-series 50 MHz clock signal
    input wire [9:0] SW;        // DE-series switches
    input wire [3:0] KEY;       // DE-series pushbuttons
    output wire [9:0] LEDR;     // DE-series LEDs   

    Counter U1 (KEY[0], CLOCK_50, LEDR);

endmodule

